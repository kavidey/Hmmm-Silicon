VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hmmm
  CLASS BLOCK ;
  FOREIGN hmmm ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1230.840 4.000 1231.440 ;
    END
  END clk
  PIN halt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 207.440 1499.000 208.040 ;
    END
  END halt
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 768.440 1499.000 769.040 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1455.240 4.000 1455.840 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 880.640 1499.000 881.240 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1118.640 4.000 1119.240 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 95.240 1499.000 95.840 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 1.000 1272.270 4.000 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 1.000 1059.750 4.000 ;
    END
  END in[15]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1496.000 1127.370 1499.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1.000 315.930 4.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 319.640 1499.000 320.240 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1496.000 914.850 1499.000 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 333.240 4.000 333.840 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 445.440 4.000 446.040 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 431.840 1499.000 432.440 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1105.040 1499.000 1105.640 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1496.000 64.770 1499.000 ;
    END
  END in[9]
  PIN oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1.000 847.230 4.000 ;
    END
  END oeb[0]
  PIN oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1441.640 1499.000 1442.240 ;
    END
  END oeb[10]
  PIN oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 1.000 1166.010 4.000 ;
    END
  END oeb[11]
  PIN oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 1496.000 277.290 1499.000 ;
    END
  END oeb[12]
  PIN oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 782.040 4.000 782.640 ;
    END
  END oeb[13]
  PIN oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 1.000 1484.790 4.000 ;
    END
  END oeb[14]
  PIN oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1496.000 596.070 1499.000 ;
    END
  END oeb[15]
  PIN oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1496.000 1233.630 1499.000 ;
    END
  END oeb[1]
  PIN oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 221.040 4.000 221.640 ;
    END
  END oeb[2]
  PIN oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1496.000 808.590 1499.000 ;
    END
  END oeb[3]
  PIN oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1.000 634.710 4.000 ;
    END
  END oeb[4]
  PIN oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 894.240 4.000 894.840 ;
    END
  END oeb[5]
  PIN oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1217.240 1499.000 1217.840 ;
    END
  END oeb[6]
  PIN oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1496.000 171.030 1499.000 ;
    END
  END oeb[7]
  PIN oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1496.000 1021.110 1499.000 ;
    END
  END oeb[8]
  PIN oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1.000 103.410 4.000 ;
    END
  END oeb[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 669.840 4.000 670.440 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1329.440 1499.000 1330.040 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1.000 528.450 4.000 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 992.840 1499.000 993.440 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 1.000 1378.530 4.000 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1496.000 702.330 1499.000 ;
    END
  END out[15]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 544.040 1499.000 544.640 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1.000 209.670 4.000 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1.000 422.190 4.000 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1006.440 4.000 1007.040 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.840 4.000 109.440 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1.000 740.970 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 1496.000 1446.150 1499.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 1496.000 1339.890 1499.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1496.000 383.550 1499.000 ;
    END
  END out[9]
  PIN pgrm_addr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1496.000 489.810 1499.000 ;
    END
  END pgrm_addr
  PIN pgrm_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1.000 953.490 4.000 ;
    END
  END pgrm_data
  PIN read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 557.640 4.000 558.240 ;
    END
  END read
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1343.040 4.000 1343.640 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  PIN write
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 656.240 1499.000 656.840 ;
    END
  END write
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 0.070 6.500 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 0.100 1495.720 64.210 1496.410 ;
        RECT 65.050 1495.720 170.470 1496.410 ;
        RECT 171.310 1495.720 276.730 1496.410 ;
        RECT 277.570 1495.720 382.990 1496.410 ;
        RECT 383.830 1495.720 489.250 1496.410 ;
        RECT 490.090 1495.720 595.510 1496.410 ;
        RECT 596.350 1495.720 701.770 1496.410 ;
        RECT 702.610 1495.720 808.030 1496.410 ;
        RECT 808.870 1495.720 914.290 1496.410 ;
        RECT 915.130 1495.720 1020.550 1496.410 ;
        RECT 1021.390 1495.720 1126.810 1496.410 ;
        RECT 1127.650 1495.720 1233.070 1496.410 ;
        RECT 1233.910 1495.720 1339.330 1496.410 ;
        RECT 1340.170 1495.720 1445.590 1496.410 ;
        RECT 1446.430 1495.720 1492.150 1496.410 ;
        RECT 0.100 4.280 1492.150 1495.720 ;
        RECT 0.650 4.000 102.850 4.280 ;
        RECT 103.690 4.000 209.110 4.280 ;
        RECT 209.950 4.000 315.370 4.280 ;
        RECT 316.210 4.000 421.630 4.280 ;
        RECT 422.470 4.000 527.890 4.280 ;
        RECT 528.730 4.000 634.150 4.280 ;
        RECT 634.990 4.000 740.410 4.280 ;
        RECT 741.250 4.000 846.670 4.280 ;
        RECT 847.510 4.000 952.930 4.280 ;
        RECT 953.770 4.000 1059.190 4.280 ;
        RECT 1060.030 4.000 1165.450 4.280 ;
        RECT 1166.290 4.000 1271.710 4.280 ;
        RECT 1272.550 4.000 1377.970 4.280 ;
        RECT 1378.810 4.000 1484.230 4.280 ;
        RECT 1485.070 4.000 1492.150 4.280 ;
      LAYER met3 ;
        RECT 4.000 1456.240 1496.000 1488.005 ;
        RECT 4.400 1454.840 1496.000 1456.240 ;
        RECT 4.000 1442.640 1496.000 1454.840 ;
        RECT 4.000 1441.240 1495.600 1442.640 ;
        RECT 4.000 1344.040 1496.000 1441.240 ;
        RECT 4.400 1342.640 1496.000 1344.040 ;
        RECT 4.000 1330.440 1496.000 1342.640 ;
        RECT 4.000 1329.040 1495.600 1330.440 ;
        RECT 4.000 1231.840 1496.000 1329.040 ;
        RECT 4.400 1230.440 1496.000 1231.840 ;
        RECT 4.000 1218.240 1496.000 1230.440 ;
        RECT 4.000 1216.840 1495.600 1218.240 ;
        RECT 4.000 1119.640 1496.000 1216.840 ;
        RECT 4.400 1118.240 1496.000 1119.640 ;
        RECT 4.000 1106.040 1496.000 1118.240 ;
        RECT 4.000 1104.640 1495.600 1106.040 ;
        RECT 4.000 1007.440 1496.000 1104.640 ;
        RECT 4.400 1006.040 1496.000 1007.440 ;
        RECT 4.000 993.840 1496.000 1006.040 ;
        RECT 4.000 992.440 1495.600 993.840 ;
        RECT 4.000 895.240 1496.000 992.440 ;
        RECT 4.400 893.840 1496.000 895.240 ;
        RECT 4.000 881.640 1496.000 893.840 ;
        RECT 4.000 880.240 1495.600 881.640 ;
        RECT 4.000 783.040 1496.000 880.240 ;
        RECT 4.400 781.640 1496.000 783.040 ;
        RECT 4.000 769.440 1496.000 781.640 ;
        RECT 4.000 768.040 1495.600 769.440 ;
        RECT 4.000 670.840 1496.000 768.040 ;
        RECT 4.400 669.440 1496.000 670.840 ;
        RECT 4.000 657.240 1496.000 669.440 ;
        RECT 4.000 655.840 1495.600 657.240 ;
        RECT 4.000 558.640 1496.000 655.840 ;
        RECT 4.400 557.240 1496.000 558.640 ;
        RECT 4.000 545.040 1496.000 557.240 ;
        RECT 4.000 543.640 1495.600 545.040 ;
        RECT 4.000 446.440 1496.000 543.640 ;
        RECT 4.400 445.040 1496.000 446.440 ;
        RECT 4.000 432.840 1496.000 445.040 ;
        RECT 4.000 431.440 1495.600 432.840 ;
        RECT 4.000 334.240 1496.000 431.440 ;
        RECT 4.400 332.840 1496.000 334.240 ;
        RECT 4.000 320.640 1496.000 332.840 ;
        RECT 4.000 319.240 1495.600 320.640 ;
        RECT 4.000 222.040 1496.000 319.240 ;
        RECT 4.400 220.640 1496.000 222.040 ;
        RECT 4.000 208.440 1496.000 220.640 ;
        RECT 4.000 207.040 1495.600 208.440 ;
        RECT 4.000 109.840 1496.000 207.040 ;
        RECT 4.400 108.440 1496.000 109.840 ;
        RECT 4.000 96.240 1496.000 108.440 ;
        RECT 4.000 94.840 1495.600 96.240 ;
        RECT 4.000 10.715 1496.000 94.840 ;
      LAYER met4 ;
        RECT 228.455 11.735 251.040 1486.305 ;
        RECT 253.440 11.735 327.840 1486.305 ;
        RECT 330.240 11.735 404.640 1486.305 ;
        RECT 407.040 11.735 481.440 1486.305 ;
        RECT 483.840 11.735 558.240 1486.305 ;
        RECT 560.640 11.735 635.040 1486.305 ;
        RECT 637.440 11.735 711.840 1486.305 ;
        RECT 714.240 11.735 788.640 1486.305 ;
        RECT 791.040 11.735 865.440 1486.305 ;
        RECT 867.840 11.735 942.240 1486.305 ;
        RECT 944.640 11.735 1019.040 1486.305 ;
        RECT 1021.440 11.735 1095.840 1486.305 ;
        RECT 1098.240 11.735 1172.640 1486.305 ;
        RECT 1175.040 11.735 1249.440 1486.305 ;
        RECT 1251.840 11.735 1284.945 1486.305 ;
  END
END hmmm
END LIBRARY

