VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hmmm
  CLASS BLOCK ;
  FOREIGN hmmm ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.000 BY 3000.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2043.440 4.000 2044.040 ;
    END
  END clk
  PIN halt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 860.240 1999.000 860.840 ;
    END
  END halt
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1791.840 1999.000 1792.440 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2417.440 4.000 2418.040 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1978.840 1999.000 1979.440 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1859.840 4.000 1860.440 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 673.240 1999.000 673.840 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 115.640 1999.000 116.240 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 1.000 1761.710 4.000 ;
    END
  END in[15]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 2996.000 1384.970 2999.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1.000 528.450 4.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1047.240 1999.000 1047.840 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 2996.000 1030.770 2999.000 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 557.640 4.000 558.240 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 741.240 4.000 741.840 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1234.240 1999.000 1234.840 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2349.440 1999.000 2350.040 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2604.440 4.000 2605.040 ;
    END
  END in[9]
  PIN oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1.000 1407.510 4.000 ;
    END
  END oeb[0]
  PIN oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2907.040 1999.000 2907.640 ;
    END
  END oeb[10]
  PIN oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 1.000 1938.810 4.000 ;
    END
  END oeb[11]
  PIN oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2975.040 4.000 2975.640 ;
    END
  END oeb[12]
  PIN oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1302.240 4.000 1302.840 ;
    END
  END oeb[13]
  PIN oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 489.640 1999.000 490.240 ;
    END
  END oeb[14]
  PIN oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 2996.000 502.690 2999.000 ;
    END
  END oeb[15]
  PIN oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 2996.000 1562.070 2999.000 ;
    END
  END oeb[1]
  PIN oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 370.640 4.000 371.240 ;
    END
  END oeb[2]
  PIN oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 2996.000 856.890 2999.000 ;
    END
  END oeb[3]
  PIN oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1.000 1056.530 4.000 ;
    END
  END oeb[4]
  PIN oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1485.840 4.000 1486.440 ;
    END
  END oeb[5]
  PIN oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2536.440 1999.000 2537.040 ;
    END
  END oeb[6]
  PIN oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2788.040 4.000 2788.640 ;
    END
  END oeb[7]
  PIN oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 2996.000 1207.870 2999.000 ;
    END
  END oeb[8]
  PIN oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1.000 174.250 4.000 ;
    END
  END oeb[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1115.240 4.000 1115.840 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2720.040 1999.000 2720.640 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1.000 879.430 4.000 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2162.440 1999.000 2163.040 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 302.640 1999.000 303.240 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 2996.000 679.790 2999.000 ;
    END
  END out[15]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1417.840 1999.000 1418.440 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 1.000 351.350 4.000 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1.000 702.330 4.000 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1672.840 4.000 1673.440 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.640 4.000 184.240 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1.000 1233.630 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 2996.000 1913.050 2999.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 2996.000 1735.950 2999.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 2996.000 151.710 2999.000 ;
    END
  END out[9]
  PIN pgrm_addr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 2996.000 328.810 2999.000 ;
    END
  END pgrm_addr
  PIN pgrm_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 1.000 1584.610 4.000 ;
    END
  END pgrm_data
  PIN read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 928.240 4.000 928.840 ;
    END
  END read
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 2230.440 4.000 2231.040 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2986.800 ;
    END
  END vssd1
  PIN write
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1604.840 1999.000 1605.440 ;
    END
  END write
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1994.100 2986.645 ;
      LAYER met1 ;
        RECT 0.070 6.500 1994.100 2986.800 ;
      LAYER met2 ;
        RECT 0.100 2995.720 151.150 2996.490 ;
        RECT 151.990 2995.720 328.250 2996.490 ;
        RECT 329.090 2995.720 502.130 2996.490 ;
        RECT 502.970 2995.720 679.230 2996.490 ;
        RECT 680.070 2995.720 856.330 2996.490 ;
        RECT 857.170 2995.720 1030.210 2996.490 ;
        RECT 1031.050 2995.720 1207.310 2996.490 ;
        RECT 1208.150 2995.720 1384.410 2996.490 ;
        RECT 1385.250 2995.720 1561.510 2996.490 ;
        RECT 1562.350 2995.720 1735.390 2996.490 ;
        RECT 1736.230 2995.720 1912.490 2996.490 ;
        RECT 1913.330 2995.720 1992.620 2996.490 ;
        RECT 0.100 4.280 1992.620 2995.720 ;
        RECT 0.650 3.670 173.690 4.280 ;
        RECT 174.530 3.670 350.790 4.280 ;
        RECT 351.630 3.670 527.890 4.280 ;
        RECT 528.730 3.670 701.770 4.280 ;
        RECT 702.610 3.670 878.870 4.280 ;
        RECT 879.710 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1233.070 4.280 ;
        RECT 1233.910 3.670 1406.950 4.280 ;
        RECT 1407.790 3.670 1584.050 4.280 ;
        RECT 1584.890 3.670 1761.150 4.280 ;
        RECT 1761.990 3.670 1938.250 4.280 ;
        RECT 1939.090 3.670 1992.620 4.280 ;
      LAYER met3 ;
        RECT 4.000 2976.040 1996.000 2986.725 ;
        RECT 4.400 2974.640 1996.000 2976.040 ;
        RECT 4.000 2908.040 1996.000 2974.640 ;
        RECT 4.000 2906.640 1995.600 2908.040 ;
        RECT 4.000 2789.040 1996.000 2906.640 ;
        RECT 4.400 2787.640 1996.000 2789.040 ;
        RECT 4.000 2721.040 1996.000 2787.640 ;
        RECT 4.000 2719.640 1995.600 2721.040 ;
        RECT 4.000 2605.440 1996.000 2719.640 ;
        RECT 4.400 2604.040 1996.000 2605.440 ;
        RECT 4.000 2537.440 1996.000 2604.040 ;
        RECT 4.000 2536.040 1995.600 2537.440 ;
        RECT 4.000 2418.440 1996.000 2536.040 ;
        RECT 4.400 2417.040 1996.000 2418.440 ;
        RECT 4.000 2350.440 1996.000 2417.040 ;
        RECT 4.000 2349.040 1995.600 2350.440 ;
        RECT 4.000 2231.440 1996.000 2349.040 ;
        RECT 4.400 2230.040 1996.000 2231.440 ;
        RECT 4.000 2163.440 1996.000 2230.040 ;
        RECT 4.000 2162.040 1995.600 2163.440 ;
        RECT 4.000 2044.440 1996.000 2162.040 ;
        RECT 4.400 2043.040 1996.000 2044.440 ;
        RECT 4.000 1979.840 1996.000 2043.040 ;
        RECT 4.000 1978.440 1995.600 1979.840 ;
        RECT 4.000 1860.840 1996.000 1978.440 ;
        RECT 4.400 1859.440 1996.000 1860.840 ;
        RECT 4.000 1792.840 1996.000 1859.440 ;
        RECT 4.000 1791.440 1995.600 1792.840 ;
        RECT 4.000 1673.840 1996.000 1791.440 ;
        RECT 4.400 1672.440 1996.000 1673.840 ;
        RECT 4.000 1605.840 1996.000 1672.440 ;
        RECT 4.000 1604.440 1995.600 1605.840 ;
        RECT 4.000 1486.840 1996.000 1604.440 ;
        RECT 4.400 1485.440 1996.000 1486.840 ;
        RECT 4.000 1418.840 1996.000 1485.440 ;
        RECT 4.000 1417.440 1995.600 1418.840 ;
        RECT 4.000 1303.240 1996.000 1417.440 ;
        RECT 4.400 1301.840 1996.000 1303.240 ;
        RECT 4.000 1235.240 1996.000 1301.840 ;
        RECT 4.000 1233.840 1995.600 1235.240 ;
        RECT 4.000 1116.240 1996.000 1233.840 ;
        RECT 4.400 1114.840 1996.000 1116.240 ;
        RECT 4.000 1048.240 1996.000 1114.840 ;
        RECT 4.000 1046.840 1995.600 1048.240 ;
        RECT 4.000 929.240 1996.000 1046.840 ;
        RECT 4.400 927.840 1996.000 929.240 ;
        RECT 4.000 861.240 1996.000 927.840 ;
        RECT 4.000 859.840 1995.600 861.240 ;
        RECT 4.000 742.240 1996.000 859.840 ;
        RECT 4.400 740.840 1996.000 742.240 ;
        RECT 4.000 674.240 1996.000 740.840 ;
        RECT 4.000 672.840 1995.600 674.240 ;
        RECT 4.000 558.640 1996.000 672.840 ;
        RECT 4.400 557.240 1996.000 558.640 ;
        RECT 4.000 490.640 1996.000 557.240 ;
        RECT 4.000 489.240 1995.600 490.640 ;
        RECT 4.000 371.640 1996.000 489.240 ;
        RECT 4.400 370.240 1996.000 371.640 ;
        RECT 4.000 303.640 1996.000 370.240 ;
        RECT 4.000 302.240 1995.600 303.640 ;
        RECT 4.000 184.640 1996.000 302.240 ;
        RECT 4.400 183.240 1996.000 184.640 ;
        RECT 4.000 116.640 1996.000 183.240 ;
        RECT 4.000 115.240 1995.600 116.640 ;
        RECT 4.000 10.715 1996.000 115.240 ;
      LAYER met4 ;
        RECT 551.375 15.135 558.240 2039.145 ;
        RECT 560.640 15.135 635.040 2039.145 ;
        RECT 637.440 15.135 711.840 2039.145 ;
        RECT 714.240 15.135 788.640 2039.145 ;
        RECT 791.040 15.135 865.440 2039.145 ;
        RECT 867.840 15.135 942.240 2039.145 ;
        RECT 944.640 15.135 1019.040 2039.145 ;
        RECT 1021.440 15.135 1095.840 2039.145 ;
        RECT 1098.240 15.135 1172.640 2039.145 ;
        RECT 1175.040 15.135 1249.440 2039.145 ;
        RECT 1251.840 15.135 1326.240 2039.145 ;
        RECT 1328.640 15.135 1403.040 2039.145 ;
        RECT 1405.440 15.135 1477.225 2039.145 ;
  END
END hmmm
END LIBRARY

