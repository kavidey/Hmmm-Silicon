magic
tech sky130A
magscale 1 2
timestamp 1673295837
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 14 1300 298816 297616
<< metal2 >>
rect 12898 299200 12954 299800
rect 34150 299200 34206 299800
rect 55402 299200 55458 299800
rect 76654 299200 76710 299800
rect 97906 299200 97962 299800
rect 119158 299200 119214 299800
rect 140410 299200 140466 299800
rect 161662 299200 161718 299800
rect 182914 299200 182970 299800
rect 204166 299200 204222 299800
rect 225418 299200 225474 299800
rect 246670 299200 246726 299800
rect 267922 299200 267978 299800
rect 289174 299200 289230 299800
rect 18 200 74 800
rect 20626 200 20682 800
rect 41878 200 41934 800
rect 63130 200 63186 800
rect 84382 200 84438 800
rect 105634 200 105690 800
rect 126886 200 126942 800
rect 148138 200 148194 800
rect 169390 200 169446 800
rect 190642 200 190698 800
rect 211894 200 211950 800
rect 233146 200 233202 800
rect 254398 200 254454 800
rect 275650 200 275706 800
rect 296902 200 296958 800
<< obsm2 >>
rect 20 299144 12842 299282
rect 13010 299144 34094 299282
rect 34262 299144 55346 299282
rect 55514 299144 76598 299282
rect 76766 299144 97850 299282
rect 98018 299144 119102 299282
rect 119270 299144 140354 299282
rect 140522 299144 161606 299282
rect 161774 299144 182858 299282
rect 183026 299144 204110 299282
rect 204278 299144 225362 299282
rect 225530 299144 246614 299282
rect 246782 299144 267866 299282
rect 268034 299144 289118 299282
rect 289286 299144 298430 299282
rect 20 856 298430 299144
rect 130 800 20570 856
rect 20738 800 41822 856
rect 41990 800 63074 856
rect 63242 800 84326 856
rect 84494 800 105578 856
rect 105746 800 126830 856
rect 126998 800 148082 856
rect 148250 800 169334 856
rect 169502 800 190586 856
rect 190754 800 211838 856
rect 212006 800 233090 856
rect 233258 800 254342 856
rect 254510 800 275594 856
rect 275762 800 296846 856
rect 297014 800 298430 856
<< metal3 >>
rect 200 291048 800 291168
rect 299200 288328 299800 288448
rect 200 268608 800 268728
rect 299200 265888 299800 266008
rect 200 246168 800 246288
rect 299200 243448 299800 243568
rect 200 223728 800 223848
rect 299200 221008 299800 221128
rect 200 201288 800 201408
rect 299200 198568 299800 198688
rect 200 178848 800 178968
rect 299200 176128 299800 176248
rect 200 156408 800 156528
rect 299200 153688 299800 153808
rect 200 133968 800 134088
rect 299200 131248 299800 131368
rect 200 111528 800 111648
rect 299200 108808 299800 108928
rect 200 89088 800 89208
rect 299200 86368 299800 86488
rect 200 66648 800 66768
rect 299200 63928 299800 64048
rect 200 44208 800 44328
rect 299200 41488 299800 41608
rect 200 21768 800 21888
rect 299200 19048 299800 19168
<< obsm3 >>
rect 800 291248 299200 297601
rect 880 290968 299200 291248
rect 800 288528 299200 290968
rect 800 288248 299120 288528
rect 800 268808 299200 288248
rect 880 268528 299200 268808
rect 800 266088 299200 268528
rect 800 265808 299120 266088
rect 800 246368 299200 265808
rect 880 246088 299200 246368
rect 800 243648 299200 246088
rect 800 243368 299120 243648
rect 800 223928 299200 243368
rect 880 223648 299200 223928
rect 800 221208 299200 223648
rect 800 220928 299120 221208
rect 800 201488 299200 220928
rect 880 201208 299200 201488
rect 800 198768 299200 201208
rect 800 198488 299120 198768
rect 800 179048 299200 198488
rect 880 178768 299200 179048
rect 800 176328 299200 178768
rect 800 176048 299120 176328
rect 800 156608 299200 176048
rect 880 156328 299200 156608
rect 800 153888 299200 156328
rect 800 153608 299120 153888
rect 800 134168 299200 153608
rect 880 133888 299200 134168
rect 800 131448 299200 133888
rect 800 131168 299120 131448
rect 800 111728 299200 131168
rect 880 111448 299200 111728
rect 800 109008 299200 111448
rect 800 108728 299120 109008
rect 800 89288 299200 108728
rect 880 89008 299200 89288
rect 800 86568 299200 89008
rect 800 86288 299120 86568
rect 800 66848 299200 86288
rect 880 66568 299200 66848
rect 800 64128 299200 66568
rect 800 63848 299120 64128
rect 800 44408 299200 63848
rect 880 44128 299200 44408
rect 800 41688 299200 44128
rect 800 41408 299120 41688
rect 800 21968 299200 41408
rect 880 21688 299200 21968
rect 800 19248 299200 21688
rect 800 18968 299120 19248
rect 800 2143 299200 18968
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 45691 2347 50208 297261
rect 50688 2347 65568 297261
rect 66048 2347 80928 297261
rect 81408 2347 96288 297261
rect 96768 2347 111648 297261
rect 112128 2347 127008 297261
rect 127488 2347 142368 297261
rect 142848 2347 157728 297261
rect 158208 2347 173088 297261
rect 173568 2347 188448 297261
rect 188928 2347 203808 297261
rect 204288 2347 219168 297261
rect 219648 2347 234528 297261
rect 235008 2347 249888 297261
rect 250368 2347 256989 297261
<< labels >>
rlabel metal3 s 200 246168 800 246288 6 clk
port 1 nsew signal input
rlabel metal3 s 299200 41488 299800 41608 6 halt
port 2 nsew signal output
rlabel metal3 s 299200 153688 299800 153808 6 in[0]
port 3 nsew signal input
rlabel metal3 s 200 291048 800 291168 6 in[10]
port 4 nsew signal input
rlabel metal3 s 299200 176128 299800 176248 6 in[11]
port 5 nsew signal input
rlabel metal3 s 200 223728 800 223848 6 in[12]
port 6 nsew signal input
rlabel metal3 s 299200 19048 299800 19168 6 in[13]
port 7 nsew signal input
rlabel metal2 s 254398 200 254454 800 6 in[14]
port 8 nsew signal input
rlabel metal2 s 211894 200 211950 800 6 in[15]
port 9 nsew signal input
rlabel metal2 s 225418 299200 225474 299800 6 in[1]
port 10 nsew signal input
rlabel metal2 s 63130 200 63186 800 6 in[2]
port 11 nsew signal input
rlabel metal3 s 299200 63928 299800 64048 6 in[3]
port 12 nsew signal input
rlabel metal2 s 182914 299200 182970 299800 6 in[4]
port 13 nsew signal input
rlabel metal3 s 200 66648 800 66768 6 in[5]
port 14 nsew signal input
rlabel metal3 s 200 89088 800 89208 6 in[6]
port 15 nsew signal input
rlabel metal3 s 299200 86368 299800 86488 6 in[7]
port 16 nsew signal input
rlabel metal3 s 299200 221008 299800 221128 6 in[8]
port 17 nsew signal input
rlabel metal2 s 12898 299200 12954 299800 6 in[9]
port 18 nsew signal input
rlabel metal2 s 169390 200 169446 800 6 oeb[0]
port 19 nsew signal output
rlabel metal3 s 299200 288328 299800 288448 6 oeb[10]
port 20 nsew signal output
rlabel metal2 s 233146 200 233202 800 6 oeb[11]
port 21 nsew signal output
rlabel metal2 s 55402 299200 55458 299800 6 oeb[12]
port 22 nsew signal output
rlabel metal3 s 200 156408 800 156528 6 oeb[13]
port 23 nsew signal output
rlabel metal2 s 296902 200 296958 800 6 oeb[14]
port 24 nsew signal output
rlabel metal2 s 119158 299200 119214 299800 6 oeb[15]
port 25 nsew signal output
rlabel metal2 s 246670 299200 246726 299800 6 oeb[1]
port 26 nsew signal output
rlabel metal3 s 200 44208 800 44328 6 oeb[2]
port 27 nsew signal output
rlabel metal2 s 161662 299200 161718 299800 6 oeb[3]
port 28 nsew signal output
rlabel metal2 s 126886 200 126942 800 6 oeb[4]
port 29 nsew signal output
rlabel metal3 s 200 178848 800 178968 6 oeb[5]
port 30 nsew signal output
rlabel metal3 s 299200 243448 299800 243568 6 oeb[6]
port 31 nsew signal output
rlabel metal2 s 34150 299200 34206 299800 6 oeb[7]
port 32 nsew signal output
rlabel metal2 s 204166 299200 204222 299800 6 oeb[8]
port 33 nsew signal output
rlabel metal2 s 20626 200 20682 800 6 oeb[9]
port 34 nsew signal output
rlabel metal2 s 18 200 74 800 6 out[0]
port 35 nsew signal output
rlabel metal3 s 200 133968 800 134088 6 out[10]
port 36 nsew signal output
rlabel metal3 s 299200 265888 299800 266008 6 out[11]
port 37 nsew signal output
rlabel metal2 s 105634 200 105690 800 6 out[12]
port 38 nsew signal output
rlabel metal3 s 299200 198568 299800 198688 6 out[13]
port 39 nsew signal output
rlabel metal2 s 275650 200 275706 800 6 out[14]
port 40 nsew signal output
rlabel metal2 s 140410 299200 140466 299800 6 out[15]
port 41 nsew signal output
rlabel metal3 s 299200 108808 299800 108928 6 out[1]
port 42 nsew signal output
rlabel metal2 s 41878 200 41934 800 6 out[2]
port 43 nsew signal output
rlabel metal2 s 84382 200 84438 800 6 out[3]
port 44 nsew signal output
rlabel metal3 s 200 201288 800 201408 6 out[4]
port 45 nsew signal output
rlabel metal3 s 200 21768 800 21888 6 out[5]
port 46 nsew signal output
rlabel metal2 s 148138 200 148194 800 6 out[6]
port 47 nsew signal output
rlabel metal2 s 289174 299200 289230 299800 6 out[7]
port 48 nsew signal output
rlabel metal2 s 267922 299200 267978 299800 6 out[8]
port 49 nsew signal output
rlabel metal2 s 76654 299200 76710 299800 6 out[9]
port 50 nsew signal output
rlabel metal2 s 97906 299200 97962 299800 6 pgrm_addr
port 51 nsew signal input
rlabel metal2 s 190642 200 190698 800 6 pgrm_data
port 52 nsew signal input
rlabel metal3 s 200 111528 800 111648 6 read
port 53 nsew signal output
rlabel metal3 s 200 268608 800 268728 6 rst
port 54 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 56 nsew ground bidirectional
rlabel metal3 s 299200 131248 299800 131368 6 write
port 57 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 112068446
string GDS_FILE /Users/kavidey/github/Hmmm-Silicon/openlane/hmmm/runs/23_01_09_11_38/results/signoff/hmmm.magic.gds
string GDS_START 1198492
<< end >>

