magic
tech sky130A
magscale 1 2
timestamp 1673602232
<< obsli1 >>
rect 1104 2159 398820 597329
<< obsm1 >>
rect 14 1300 398820 597360
<< metal2 >>
rect 30286 599200 30342 599800
rect 65706 599200 65762 599800
rect 100482 599200 100538 599800
rect 135902 599200 135958 599800
rect 171322 599200 171378 599800
rect 206098 599200 206154 599800
rect 241518 599200 241574 599800
rect 276938 599200 276994 599800
rect 312358 599200 312414 599800
rect 347134 599200 347190 599800
rect 382554 599200 382610 599800
rect 18 200 74 800
rect 34794 200 34850 800
rect 70214 200 70270 800
rect 105634 200 105690 800
rect 140410 200 140466 800
rect 175830 200 175886 800
rect 211250 200 211306 800
rect 246670 200 246726 800
rect 281446 200 281502 800
rect 316866 200 316922 800
rect 352286 200 352342 800
rect 387706 200 387762 800
<< obsm2 >>
rect 20 599144 30230 599298
rect 30398 599144 65650 599298
rect 65818 599144 100426 599298
rect 100594 599144 135846 599298
rect 136014 599144 171266 599298
rect 171434 599144 206042 599298
rect 206210 599144 241462 599298
rect 241630 599144 276882 599298
rect 277050 599144 312302 599298
rect 312470 599144 347078 599298
rect 347246 599144 382498 599298
rect 382666 599144 398434 599298
rect 20 856 398434 599144
rect 130 800 34738 856
rect 34906 800 70158 856
rect 70326 800 105578 856
rect 105746 800 140354 856
rect 140522 800 175774 856
rect 175942 800 211194 856
rect 211362 800 246614 856
rect 246782 800 281390 856
rect 281558 800 316810 856
rect 316978 800 352230 856
rect 352398 800 387650 856
rect 387818 800 398434 856
<< metal3 >>
rect 200 595008 800 595128
rect 399200 581408 399800 581528
rect 200 557608 800 557728
rect 399200 544008 399800 544128
rect 200 520888 800 521008
rect 399200 507288 399800 507408
rect 200 483488 800 483608
rect 399200 469888 399800 470008
rect 200 446088 800 446208
rect 399200 432488 399800 432608
rect 200 408688 800 408808
rect 399200 395768 399800 395888
rect 200 371968 800 372088
rect 399200 358368 399800 358488
rect 200 334568 800 334688
rect 399200 320968 399800 321088
rect 200 297168 800 297288
rect 399200 283568 399800 283688
rect 200 260448 800 260568
rect 399200 246848 399800 246968
rect 200 223048 800 223168
rect 399200 209448 399800 209568
rect 200 185648 800 185768
rect 399200 172048 399800 172168
rect 200 148248 800 148368
rect 399200 134648 399800 134768
rect 200 111528 800 111648
rect 399200 97928 399800 98048
rect 200 74128 800 74248
rect 399200 60528 399800 60648
rect 200 36728 800 36848
rect 399200 23128 399800 23248
<< obsm3 >>
rect 800 595208 399200 597345
rect 880 594928 399200 595208
rect 800 581608 399200 594928
rect 800 581328 399120 581608
rect 800 557808 399200 581328
rect 880 557528 399200 557808
rect 800 544208 399200 557528
rect 800 543928 399120 544208
rect 800 521088 399200 543928
rect 880 520808 399200 521088
rect 800 507488 399200 520808
rect 800 507208 399120 507488
rect 800 483688 399200 507208
rect 880 483408 399200 483688
rect 800 470088 399200 483408
rect 800 469808 399120 470088
rect 800 446288 399200 469808
rect 880 446008 399200 446288
rect 800 432688 399200 446008
rect 800 432408 399120 432688
rect 800 408888 399200 432408
rect 880 408608 399200 408888
rect 800 395968 399200 408608
rect 800 395688 399120 395968
rect 800 372168 399200 395688
rect 880 371888 399200 372168
rect 800 358568 399200 371888
rect 800 358288 399120 358568
rect 800 334768 399200 358288
rect 880 334488 399200 334768
rect 800 321168 399200 334488
rect 800 320888 399120 321168
rect 800 297368 399200 320888
rect 880 297088 399200 297368
rect 800 283768 399200 297088
rect 800 283488 399120 283768
rect 800 260648 399200 283488
rect 880 260368 399200 260648
rect 800 247048 399200 260368
rect 800 246768 399120 247048
rect 800 223248 399200 246768
rect 880 222968 399200 223248
rect 800 209648 399200 222968
rect 800 209368 399120 209648
rect 800 185848 399200 209368
rect 880 185568 399200 185848
rect 800 172248 399200 185568
rect 800 171968 399120 172248
rect 800 148448 399200 171968
rect 880 148168 399200 148448
rect 800 134848 399200 148168
rect 800 134568 399120 134848
rect 800 111728 399200 134568
rect 880 111448 399200 111728
rect 800 98128 399200 111448
rect 800 97848 399120 98128
rect 800 74328 399200 97848
rect 880 74048 399200 74328
rect 800 60728 399200 74048
rect 800 60448 399120 60728
rect 800 36928 399200 60448
rect 880 36648 399200 36928
rect 800 23328 399200 36648
rect 800 23048 399120 23328
rect 800 2143 399200 23048
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
rect 111728 2128 112048 597360
rect 127088 2128 127408 597360
rect 142448 2128 142768 597360
rect 157808 2128 158128 597360
rect 173168 2128 173488 597360
rect 188528 2128 188848 597360
rect 203888 2128 204208 597360
rect 219248 2128 219568 597360
rect 234608 2128 234928 597360
rect 249968 2128 250288 597360
rect 265328 2128 265648 597360
rect 280688 2128 281008 597360
rect 296048 2128 296368 597360
rect 311408 2128 311728 597360
rect 326768 2128 327088 597360
rect 342128 2128 342448 597360
rect 357488 2128 357808 597360
rect 372848 2128 373168 597360
rect 388208 2128 388528 597360
<< obsm4 >>
rect 112667 81363 127008 469301
rect 127488 81363 142368 469301
rect 142848 81363 157728 469301
rect 158208 81363 173088 469301
rect 173568 81363 188448 469301
rect 188928 81363 203808 469301
rect 204288 81363 219168 469301
rect 219648 81363 234528 469301
rect 235008 81363 249888 469301
rect 250368 81363 265248 469301
rect 265728 81363 280608 469301
rect 281088 81363 291029 469301
<< labels >>
rlabel metal3 s 200 408688 800 408808 6 clk
port 1 nsew signal input
rlabel metal3 s 399200 172048 399800 172168 6 halt
port 2 nsew signal output
rlabel metal3 s 399200 358368 399800 358488 6 in[0]
port 3 nsew signal input
rlabel metal3 s 200 483488 800 483608 6 in[10]
port 4 nsew signal input
rlabel metal3 s 399200 395768 399800 395888 6 in[11]
port 5 nsew signal input
rlabel metal3 s 200 371968 800 372088 6 in[12]
port 6 nsew signal input
rlabel metal3 s 399200 134648 399800 134768 6 in[13]
port 7 nsew signal input
rlabel metal3 s 399200 23128 399800 23248 6 in[14]
port 8 nsew signal input
rlabel metal2 s 352286 200 352342 800 6 in[15]
port 9 nsew signal input
rlabel metal2 s 276938 599200 276994 599800 6 in[1]
port 10 nsew signal input
rlabel metal2 s 105634 200 105690 800 6 in[2]
port 11 nsew signal input
rlabel metal3 s 399200 209448 399800 209568 6 in[3]
port 12 nsew signal input
rlabel metal2 s 206098 599200 206154 599800 6 in[4]
port 13 nsew signal input
rlabel metal3 s 200 111528 800 111648 6 in[5]
port 14 nsew signal input
rlabel metal3 s 200 148248 800 148368 6 in[6]
port 15 nsew signal input
rlabel metal3 s 399200 246848 399800 246968 6 in[7]
port 16 nsew signal input
rlabel metal3 s 399200 469888 399800 470008 6 in[8]
port 17 nsew signal input
rlabel metal3 s 200 520888 800 521008 6 in[9]
port 18 nsew signal input
rlabel metal2 s 281446 200 281502 800 6 oeb[0]
port 19 nsew signal output
rlabel metal3 s 399200 581408 399800 581528 6 oeb[10]
port 20 nsew signal output
rlabel metal2 s 387706 200 387762 800 6 oeb[11]
port 21 nsew signal output
rlabel metal3 s 200 595008 800 595128 6 oeb[12]
port 22 nsew signal output
rlabel metal3 s 200 260448 800 260568 6 oeb[13]
port 23 nsew signal output
rlabel metal3 s 399200 97928 399800 98048 6 oeb[14]
port 24 nsew signal output
rlabel metal2 s 100482 599200 100538 599800 6 oeb[15]
port 25 nsew signal output
rlabel metal2 s 312358 599200 312414 599800 6 oeb[1]
port 26 nsew signal output
rlabel metal3 s 200 74128 800 74248 6 oeb[2]
port 27 nsew signal output
rlabel metal2 s 171322 599200 171378 599800 6 oeb[3]
port 28 nsew signal output
rlabel metal2 s 211250 200 211306 800 6 oeb[4]
port 29 nsew signal output
rlabel metal3 s 200 297168 800 297288 6 oeb[5]
port 30 nsew signal output
rlabel metal3 s 399200 507288 399800 507408 6 oeb[6]
port 31 nsew signal output
rlabel metal3 s 200 557608 800 557728 6 oeb[7]
port 32 nsew signal output
rlabel metal2 s 241518 599200 241574 599800 6 oeb[8]
port 33 nsew signal output
rlabel metal2 s 34794 200 34850 800 6 oeb[9]
port 34 nsew signal output
rlabel metal2 s 18 200 74 800 6 out[0]
port 35 nsew signal output
rlabel metal3 s 200 223048 800 223168 6 out[10]
port 36 nsew signal output
rlabel metal3 s 399200 544008 399800 544128 6 out[11]
port 37 nsew signal output
rlabel metal2 s 175830 200 175886 800 6 out[12]
port 38 nsew signal output
rlabel metal3 s 399200 432488 399800 432608 6 out[13]
port 39 nsew signal output
rlabel metal3 s 399200 60528 399800 60648 6 out[14]
port 40 nsew signal output
rlabel metal2 s 135902 599200 135958 599800 6 out[15]
port 41 nsew signal output
rlabel metal3 s 399200 283568 399800 283688 6 out[1]
port 42 nsew signal output
rlabel metal2 s 70214 200 70270 800 6 out[2]
port 43 nsew signal output
rlabel metal2 s 140410 200 140466 800 6 out[3]
port 44 nsew signal output
rlabel metal3 s 200 334568 800 334688 6 out[4]
port 45 nsew signal output
rlabel metal3 s 200 36728 800 36848 6 out[5]
port 46 nsew signal output
rlabel metal2 s 246670 200 246726 800 6 out[6]
port 47 nsew signal output
rlabel metal2 s 382554 599200 382610 599800 6 out[7]
port 48 nsew signal output
rlabel metal2 s 347134 599200 347190 599800 6 out[8]
port 49 nsew signal output
rlabel metal2 s 30286 599200 30342 599800 6 out[9]
port 50 nsew signal output
rlabel metal2 s 65706 599200 65762 599800 6 pgrm_addr
port 51 nsew signal input
rlabel metal2 s 316866 200 316922 800 6 pgrm_data
port 52 nsew signal input
rlabel metal3 s 200 185648 800 185768 6 read
port 53 nsew signal output
rlabel metal3 s 200 446088 800 446208 6 rst
port 54 nsew signal input
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 597360 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 597360 6 vssd1
port 56 nsew ground bidirectional
rlabel metal3 s 399200 320968 399800 321088 6 write
port 57 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 400000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 157455058
string GDS_FILE /Users/kavidey/github/Hmmm-Silicon/openlane/hmmm/runs/23_01_13_01_02/results/signoff/hmmm.magic.gds
string GDS_START 1481550
<< end >>

